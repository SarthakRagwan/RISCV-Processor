module ALU_Decoder(ALUOp,op5,funct3,funct7,ALUControl);

    input funct7,op5;
    input [1:0]ALUOp;
    input [2:0]funct3;
    output [2:0]ALUControl;

    wire [1:0] concate={op5,funct7};

    assign ALUControl = (ALUOp == 2'b00) ? 3'b000 :
                        ((ALUOp == 2'b01) && (funct3 == 3'b000)) ? 3'b100 :
                        ((ALUOp == 2'b01) && (funct3 == 3'b001)) ? 3'b101 :
                        ((ALUOp == 2'b01) && (funct3 == 3'b100)) ? 3'b110 :
                        ((ALUOp == 2'b01) && (funct3 == 3'b101)) ? 3'b111 :

                        ((ALUOp == 2'b10) && (funct3 == 3'b010)) ? 3'b101 : 
                        ((ALUOp == 2'b10) && (funct3 == 3'b110)) ? 3'b011 : 
                        ((ALUOp == 2'b10) && (funct3 == 3'b111)) ? 3'b010 : 
                        ((ALUOp == 2'b11) && (funct3 == 3'b000)) ? 3'b000 :
                        ((ALUOp == 2'b11) && (funct3 == 3'b110)) ? 3'b011 :
                        ((ALUOp == 2'b11) && (funct3 == 3'b111)) ? 3'b010 :
                        ((ALUOp == 2'b10) && (funct3 == 3'b000) && (concate == 2'b11)) ? 3'b001 : 
                        ((ALUOp == 2'b10) && (funct3 == 3'b000) && (concate != 2'b11)) ? 3'b000 :
                                                                                       3'b000; 
endmodule