`include "PC.v"
`include "Instruction_Memory.v"
`include "Register_files.v"
`include "Sign_Extend.v"
`include "ALU.v"
`include "Control_Unit_Top.v"
`include "Data_Mem.v"
`include "PC_Adder.v"
`include "Mux.v"
module Single_Cycle_Top(clk,rst);
    
    input clk,rst;

    wire [31:0] PC_Top,RD_Instr_Top,RD1_TOP,Imm_Ext_Top,ALU_Result_Top,Read_Data_Top,PCPlus4_Top,RD2_TOP,SrcB_Top,Result_Top,PC_Target_Top,PC_Next_Top;
    wire [2:0] ALU_Control_Top;
    wire Reg_Write_Top,MemWrite_Top,ALUSrc_Top,ResultSrc_Top,Branch_Top;
    wire [1:0] ImmSrc_Top;
    wire branchSel;
    assign branchSel=Branch_Top & ALU_Result_Top[0];
    
    //PC: updates on each rising clock edge with PC_Next value depending on if branching took place or not
    PC_Module PC(
        .clk(clk),
        .rst(rst),
        .PC(PC_Top),
        .PC_Next(PC_Next_Top)
    );

    //PCNext: Generate next instruction address if no branching happens
    PC_Adder PC_Adder(
        .a(PC_Top),
        .b(32'd4),
        .c(PCPlus4_Top)
    );

    //PCNext: Generate next instruction address if branching happens
    PC_Adder PC_Banching(
                .a(PC_Top),
                .b(Imm_Ext_Top),
                .c(PC_Target_Top)
        );
    //Choose one of PCNext depend on branch&ALU_Result_Top[0]
    Mux Branchin_Mux(
                .a(PCPlus4_Top),
                .b(PC_Target_Top),
                .s(branchSel),
                .c(PC_Next_Top)
        );

    //Read instruction from IR with help of PC
    Instruction_Memory Instruction_Memory(
        .A(PC_Top),
        .rst(rst),
        .RD(RD_Instr_Top)
    );


    //Read and write data from/in registers corrsponding to input addresses 
    //Note: what need to be written is specified by WD3.
    //Where to write is specified by A3. 
    //When to write is specified by WE3.
    //From where to read is specified by A1/A2
    //Read data is found on RD1/Rd2

    //A1->RD1 and (A3,WD3,WE3) are used in I type instruction
    //A1->RD1 and A2->RD2 are used in S type intruction
    //A1->RD1, A2->RD2 and (A3,WD3,WE3) are used in R type instruction
    //A1->RD1 is used in B type instruction
    Reg_file Reg_file(
        .clk(clk),
        .rst(rst),
        .A1(RD_Instr_Top[19:15]),
        .A2(RD_Instr_Top[24:20]),
        .A3(RD_Instr_Top[11:7]),
        .WD3(Result_Top),
        .WE3(Reg_Write_Top),
        .RD1(RD1_TOP),
        .RD2(RD2_TOP)
    );
    
    //Sign extension of Imm value as per I type instruction when ImmSrc=00
    //Sign extension of Imm value as per S type instruction when ImmSrc=01
    //Sign extension of Imm value as per B type instruction when ImmSrc=10
    //No Imm field for R type at all
    Sign_Extend Sign_Extend(
        .In(RD_Instr_Top), 
        .Imm_Ext(Imm_Ext_Top),
        .ImmSrc(ImmSrc_Top)
    );


    //Controlled by ALUSrc
    //Choose ImmExt for I,S,B type instruction(ALUSrc=1)
    //Choose (A2->RD2) for R type instruction(ALUSrc=0) 
    Mux Mux_Register_to_ALU(
                            .a(RD2_TOP),
                            .b(Imm_Ext_Top),
                            .s(ALUSrc_Top),
                            .c(SrcB_Top)
    );

    //ALU operation according to ALUControl generated by control unit corresponding to opcode,f3 and f7
    //f7 is for only R type instruction
    ALU ALU(
        .A(RD1_TOP),
        .B(SrcB_Top),
        .Result(ALU_Result_Top),
        .ALUControl(ALU_Control_Top),
        .OverFlow(),
        .Carry(),
        .Zero(),
        .Negative()
    );

    //Generate many control signals corresponding to opcode and also generate ALUControl with the help of Table.
    Control_Unit_Top Control_Unit_Top(
        .Op(RD_Instr_Top[6:0]),
        .RegWrite(Reg_Write_Top),
        .ImmSrc(ImmSrc_Top),
        .ALUSrc(ALUSrc_Top),
        .MemWrite(MemWrite_Top),
        .ResultSrc(ResultSrc_Top),
        .Branch(Branch_Top),
        .funct3(RD_Instr_Top[14:12]),
        .funct7(RD_Instr_Top[31:25]),
        .ALUControl(ALU_Control_Top)
    );

    //when WE is high => Write the WD to address A 
    //when WE is low => Read the data from address A to RD.
    Data_Memory Data_Memory(
        .A(ALU_Result_Top),
        .WD(RD2_TOP),
        .clk(clk),
        .rst(rst),
        .WE(MemWrite_Top),
        .RD(Read_Data_Top)
    );

    //Any instruction which need not to read/write in/from data memory,it surpasses data memory through this mux controlled by ResultSrc
    Mux Mux_DataMemory_to_Register(
                            .a(ALU_Result_Top),
                            .b(Read_Data_Top),
                            .s(ResultSrc_Top),
                            .c(Result_Top)
    );
endmodule